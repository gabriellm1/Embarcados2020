
module niosLab2 (
	clk_clk,
	motor_name,
	reset_reset_n);	

	input		clk_clk;
	output	[3:0]	motor_name;
	input		reset_reset_n;
endmodule
